module nesConsle();

endmodule
