module nesConsle();

endmodule

